-------------------------------------------------------------------------------
--
-- Synthesizable model of TI's TMS9918A, TMS9928A, TMS9929A.
--
-- $Id: vdp18_clk_gen-c.vhd,v 1.5 2006/06/18 10:47:01 arnim Exp $
--
-------------------------------------------------------------------------------

configuration vdp18_clk_gen_rtl_c0 of vdp18_clk_gen is

    for rtl
    end for;
  
  end vdp18_clk_gen_rtl_c0;